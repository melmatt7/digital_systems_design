Keyboard_Control(//inputs
					  clk, kbd_data_ready, 
					  //outputs
					  direction, reset, read_signal
					  );

	inputs clk;
	
	outputs;