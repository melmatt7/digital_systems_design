`default_nettype none
module Flash_Address_Control (//input
										clk, start, read, waitRequest, dataValid
										//output 
										complete);